package pkg;
  import uvm_pkg::*;

    parameter int G_SYS_CLK = 40000000;
    parameter int G_BAUD = 256000;
    parameter int G_OVERSAMPLE = 16;
    parameter int G_WORD_WIDTH = 8;
    parameter bit G_PARITY_TYPE = 1'b1;

  
endpackage : pkg