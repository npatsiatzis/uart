package testbench_pkg;
  import uvm_pkg::*;

  `include "sequence_item.sv"
  `include "sequence.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "monitor_out.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "test.sv"

//   parameter int G_DATA_WIDTH = 6;
  
endpackage : testbench_pkg